module nor_gate_1bit(
	 output result,
    input A,
    input B
    
);
    nor nor_gate(result, A, B);
endmodule
