module and_gate_1bit(
	 output result,
    input A,
    input B
    
);
    and and_gate(result, A, B);
endmodule
